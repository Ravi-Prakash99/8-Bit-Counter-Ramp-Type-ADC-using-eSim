// Code your design here
module ravi_an(out,in_a,in_b);
  output out;
  input in_a,in_b;
  assign out = in_a && in_b ;
  
endmodule