* C:\Users\lenovo\eSim-Workspace\RAVI_ADC\RAVI_ADC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/9/2022 11:55:36 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U1-Pad3_ Net-_U10-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ ravi_counter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ ravi_an		
X2  Net-_X2-Pad1_ Net-_X2-Pad1_ GND GND GND out0 out1 out2 out3 out4 out5 out6 out7 dac_out GND avsddac_3v3_sky130_v2		
U9  Net-_U5-Pad10_ Net-_U5-Pad9_ Net-_U5-Pad8_ Net-_U5-Pad7_ Net-_U5-Pad6_ Net-_U5-Pad5_ Net-_U5-Pad4_ Net-_U5-Pad3_ out0 out1 out2 out3 out4 out5 out6 out7 dac_bridge_8		
v5  Net-_X2-Pad1_ GND DC		
U4  comp_out1 Net-_U1-Pad1_ adc_bridge_1		
v1  Net-_X1-Pad4_ GND DC		
v2  Net-_X1-Pad1_ GND DC		
v3  clk GND pulse		
U6  clk Net-_U1-Pad2_ adc_bridge_1		
U7  dac_out plot_v1		
scmode1  SKY130mode		
U3  clk plot_v1		
U2  comp_out1 plot_v1		
X1  Net-_X1-Pad1_ GND dac_out Net-_X1-Pad4_ comp_out1 rropamp31		
v4  reset GND pulse		
U8  reset plot_v1		
U10  reset Net-_U10-Pad2_ adc_bridge_1		
U15  out0 plot_v1		
U14  out1 plot_v1		
U13  out2 plot_v1		
U12  out3 plot_v1		
U11  out4 plot_v1		
U16  out5 plot_v1		
U17  out6 plot_v1		
U18  out7 plot_v1		

.end
